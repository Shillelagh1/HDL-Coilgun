module cg_top(

);

endmodule